// Listing 4.15
// This module come from our laboratorys
module disp_hex_mux
   (
    input wire clk, reset,
    input wire [3:0] hex3, hex2, hex1, hex0,  // hex digits
    input wire [3:0] dp_in,             // 4 decimal points
    output reg [3:0] an,  // enable 1-out-of-4 asserted low
    output reg [7:0] sseg // led segments
   );

   // constant declaration
   localparam N = 18;
   // internal signal declaration
   reg [N-1:0] q_reg;
   wire [N-1:0] q_next;
   reg [3:0] hex_in, hex0_nxt,hex1_nxt,hex2_nxt,hex3_nxt;
   reg dp;

   // N-bit counter
   // register
   always @(posedge clk, posedge reset)
      if (reset) begin
         q_reg <= 0;
         hex0_nxt <= 0;
         hex1_nxt <= 0;
         hex2_nxt <= 0;
         hex3_nxt <= 0;
       end
      else begin
         q_reg <= q_next;
         hex0_nxt <= hex0;
         hex1_nxt <= hex1;
         hex2_nxt <= hex2;
         hex3_nxt <= hex3;
      end

   // next-state logic
   assign q_next = q_reg + 1;

   // 2 MSBs of counter to control 4-to-1 multiplexing
   // and to generate active-low enable signal
   always @*
      case (q_reg[N-1:N-2])
         2'b00:
            begin
               an =  4'b1110;
               hex_in = hex0_nxt;
               dp = dp_in[0];
            end
         2'b01:
            begin
               an =  4'b1101;
               hex_in = hex1_nxt;
               dp = dp_in[1];
            end
         2'b10:
            begin
               an =  4'b1011;
               hex_in = hex2_nxt;
               dp = dp_in[2];
            end
         default:
            begin
               an =  4'b0111;
               hex_in = hex3_nxt;
               dp = dp_in[3];
            end
       endcase

   // hex to seven-segment led display
   always @*
   begin
      case(hex_in)
        4'h0: sseg[6:0] = 7'b1000000;
        4'h1: sseg[6:0]= 7'b1111001;
        4'h2: sseg[6:0] = 7'b0100100;
        4'h3: sseg[6:0] = 7'b0110000;
        4'h4: sseg[6:0] = 7'b0011001;
        4'h5: sseg[6:0] = 7'b0010010;
        4'h6: sseg[6:0] = 7'b0000010;
        4'h7: sseg[6:0] = 7'b1111000;
        4'h8: sseg[6:0] = 7'b0000000;
        4'h9: sseg[6:0] = 7'b0010000;
        4'ha: sseg[6:0] = 7'b0001000;
        4'hb: sseg[6:0] = 7'b0000011;
        4'hc: sseg[6:0] = 7'b1000110;
        4'hd: sseg[6:0] = 7'b0100001;
        4'he: sseg[6:0] = 7'b0000110;
        default: sseg[6:0] = 7'b0001110;  //4'hf
     endcase
     
     sseg[7] = dp;
   end

endmodule